`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:00:02 05/20/2015 
// Design Name: 
// Module Name:    SW7SegDisplayDriver 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SW7SegDisplayDriver(
CAT        , //Output to cathodes
ANO      , //Output to anodes
CLK         ,//Clock Input
CLEAR,  // Reset input
HOLD, //Hold input

    );
//------Output Ports-------
output[7:0]CAT;
output[3:0]ANO;
 
//------Input Ports--------
input CLK, CLEAR, HOLD;
 
//-----Internal Variables-----
reg[23:0]clkdiv;
reg[23:0]cathode;
 
reg[7:0]cat0;
reg[7:0]cat1;
reg[7:0]cat2;
reg[7:0]cat3;
 
reg[13:0]refclk;
reg[3:0]anode;
 
reg[3:0]ones;
reg[3:0]tens;
reg[3:0]hundreds;
 
reg onescnt;
reg tenscnt;
reg hundredscnt;
 
reg onesmaxcnt_en;
reg tensmaxcnt_en;
reg hundredsmaxcnt_en;
 
reg onesmaxcnt;
reg tensmaxcnt;
reg hundredsmaxcnt;
 
//---- internal signals
wire hold_in;
wire reset;
wire sysclk;

//Digital Clock Manager Module - Generated by ISE  
DCM_INCLKtoSYSCLK timebase_dcm ( .CLK_IN1(CLK), // Clock input (100MHz)
                                 .CLK_OUT1(sysclk) ); // Clock 0ut (11.538MHz)   
 
 
//------Code Starts Here-------
 
assign CAT = cathode;
assign ANO = anode;
assign reset = !CLEAR;
assign hold_in = HOLD;
 
//------- Base clkdiv - 100 Msec
always @(posedge sysclk)
 if (reset) begin
   clkdiv <= 24'b0 ;
 end
 else /// hold
 if (hold_in) begin
   clkdiv <= clkdiv;
   end /// end hold
 else
 if (clkdiv [23:20] == 4'b1010) begin // Terminal Count
  clkdiv <= 24'b0;
 end
 else begin
  clkdiv <= clkdiv + 1;
 end
 
//------- Refresh clkdiv 2KHz (500 uSec)
always @(posedge sysclk)
 if (reset) begin
  refclk <= 13'b0;
 end
 else
 begin
  refclk <= refclk + 1;
 end
 
//------- ones max count enable
always @(posedge sysclk)
 if (reset) begin
  onescnt <= 1'b0;
 end
 else
 begin
   onescnt <= onesmaxcnt;
   onesmaxcnt_en <= (onesmaxcnt & !onescnt);
 end
 
//------- tens max count enable
always @(posedge sysclk)
 if (reset) begin
  tenscnt <= 1'b0;
 end
 else
 begin
  tenscnt <= tensmaxcnt;
  tensmaxcnt_en <= (tensmaxcnt & !tenscnt);
 end
 
//------- hundreds max count enable
always @(posedge sysclk)
 if (reset) begin
  hundredscnt <= 1'b0;
 end
 else
 begin
  hundredscnt <= hundredsmaxcnt;
  hundredsmaxcnt_en <= (hundredsmaxcnt & !hundredscnt);
 end
 
//------- ones count
always @(posedge sysclk)
 if (reset) begin
  ones <= 4'b0000;
 end
 else
 if (onesmaxcnt_en == 1'b1) begin
   ones <= ones + 1;
 end
 else if (ones[3:0] == 4'b1010) begin
   ones <= 4'b0000;
 end
 
//------- tens count
always @(posedge sysclk)
 if (reset) begin
  tens <= 4'b0000;
 end
 else
 if (tensmaxcnt_en == 1'b1) begin
   tens <= tens + 1;
  end
  else if (tens[3:0] == 4'b1010) begin
   tens <= 4'b0000;
  end
 
//------- hundreds count
always @(posedge sysclk)
 if (reset) begin
  hundreds <= 4'b0000;
 end
 else
 if (hundredsmaxcnt_en == 1'b1) begin
  hundreds <= hundreds + 1;
 end
 else 
 if (hundreds[3:0] == 4'b1010) begin
  hundreds <= 4'b0000;
 end
 
// ----- mSec Base count ------
 
always@(posedge sysclk)
 if (reset) begin
  cat0 <= 8'b11000000;
  onesmaxcnt <= 1'b0;
 end
 else
 if(clkdiv [23:20] == 4'b0000) begin
  cat0 <= 8'b11000000;//0
  onesmaxcnt <= 1'b0;
 end
 else
 if (clkdiv [23:20] == 4'b0001) begin
  cat0 <= 8'b11111001;//1
 end
 else
 if (clkdiv [23:20] == 4'b0010) begin
   cat0 <= 8'b10100100;//2
 end
 else
 if (clkdiv [23:20] == 4'b0011) begin
  cat0 <= 8'b10110000;//3
 end
 else
 if (clkdiv [23:20] == 4'b0100) begin
  cat0 <= 8'b10011001;//4
 end
 else
 if (clkdiv [23:20] == 4'b0101) begin
  cat0 <= 8'b10010010;//5
 end
 else
 if (clkdiv [23:20] == 4'b0110) begin
  cat0 <= 8'b10000010;//6
 end
 else
 if (clkdiv [23:20] == 4'b0111) begin
  cat0 <= 8'b11111000;//7
 end
 else
 if (clkdiv [23:20] == 4'b1000) begin
  cat0 <= 8'b10000000;//8
 end
 else
 if (clkdiv [23:20] == 4'b1001) begin
  cat0 <= 8'b10011000;//9
 end
 else
 if (clkdiv [23:20] == 4'b1010) begin
  onesmaxcnt <= 1'b1;
 end
             
// ----- Sec count ------
always@(posedge sysclk)
 if (reset) begin
  cat1 <= 8'b11000000;
  tensmaxcnt <= 1'b0;
 end
 else
 if(ones [3:0] == 4'b0000) begin
  cat1 <= 8'b01000000;//0
  tensmaxcnt <= 1'b0;
 end
 else
 if (ones [3:0] == 4'b0001) begin
  cat1 <= 8'b01111001;//1
 end
 else
 if (ones [3:0] == 4'b0010) begin
  cat1 <= 8'b00100100;//2
 end
 else
 if (ones [3:0] == 4'b0011) begin
  cat1 <= 8'b00110000;//3
 end
 else
 if (ones [3:0] == 4'b0100) begin
  cat1 <= 8'b00011001;//4
 end
 else
 if (ones [3:0] == 4'b0101) begin
  cat1 <= 8'b00010010;//5
 end
 else
 if (ones [3:0] == 4'b0110) begin
  cat1 <= 8'b00000010;//6
 end
 else
 if (ones [3:0] == 4'b0111) begin
  cat1 <= 8'b01111000;//7
 end
 else
 if (ones [3:0] == 4'b1000) begin
  cat1 <= 8'b00000000;//8
 end
 else
 if (ones [3:0] == 4'b1001) begin
  cat1 <= 8'b00011000;//9
 end
 else
 if (ones [3:0] == 4'b1010) begin
  tensmaxcnt <= 1'b1;
 end
 
// ----- tens count ------
 
always@(posedge sysclk)
 if (reset) begin
  cat2 <= 8'b11000000;
  hundredsmaxcnt <= 1'b0;
 end
 else
 if(tens [3:0] == 4'b0000) begin
  cat2 <= 8'b11000000;//0
  hundredsmaxcnt <= 1'b0;
 end
 else
 if (tens [3:0] == 4'b0001) begin
  cat2 <= 8'b11111001;//1
 end
 else
 if (tens [3:0] == 4'b0010) begin
  cat2 <= 8'b10100100;//2
 end
 else
 if (tens [3:0] == 4'b0011) begin
  cat2 <= 8'b10110000;//3
 end
 else
 if (tens [3:0] == 4'b0100) begin
  cat2 <= 8'b10011001;//4
 end
 else
 if (tens [3:0] == 4'b0101) begin
  cat2 <= 8'b10010010;//5
 end
 else
 if (tens [3:0] == 4'b0110) begin
  cat2 <= 8'b10000010;//6
 end
 else
 if (tens [3:0] == 4'b0111) begin
  cat2 <= 8'b11111000;//7
 end
 else
 if (tens [3:0] == 4'b1000) begin
  cat2 <= 8'b10000000;//8
 end
 else
 if (tens [3:0] == 4'b1001) begin
  cat2 <= 8'b10011000;//9
 end
 else
 if (tens [3:0] == 4'b1010) begin
  hundredsmaxcnt <= 1'b1;
 end
// ----- hundreds count ------
 
always@(posedge sysclk)
 if (reset) begin
  cat3 <= 8'b11000000;
 end
 else
 if(hundreds [3:0] == 4'b0000) begin
  cat3 <= 8'b11000000;//0
 end
 else
 if (hundreds [3:0] == 4'b0001) begin
  cat3 <= 8'b11111001;//1
 end
 else
 if (hundreds [3:0] == 4'b0010) begin
  cat3 <= 8'b10100100;//2
 end
 else
 if (hundreds [3:0] == 4'b0011) begin
  cat3 <= 8'b10110000;//3
 end
 else
 if (hundreds [3:0] == 4'b0100) begin
  cat3 <= 8'b10011001;//4
 end
 else
 if (hundreds [3:0] == 4'b0101) begin
  cat3 <= 8'b10010010;//5
 end
 else
 if (hundreds [3:0] == 4'b0110) begin
  cat3 <= 8'b10000010;//6
 end
 else
 if (hundreds [3:0] == 4'b0111) begin
  cat3 <= 8'b11111000;//7
 end
 else
 if (hundreds [3:0] == 4'b1000) begin
  cat3 <= 8'b10000000;//8
 end
 else
 if (hundreds [3:0] == 4'b1001) begin
  cat3 <= 8'b10011000;//9
 end               
               
// ----- Anode Refresh/Cathode Mux ------
always@(posedge sysclk)
 if (reset) begin
  anode <= 4'B0000;
  cathode <= 8'b11000000;
 end
 else
 if(refclk [12:11] == 2'b00) begin
  anode <=4'b0001;
  cathode <= cat0;
 end
 else
 if(refclk [12:11] == 2'b01) begin
  anode <=4'b0010;
  cathode <= cat1;
 end
 else
 if(refclk [12:11] == 2'b10) begin
  anode <=4'b0100;
  cathode <= cat2;
 end
 else
 if(refclk [12:11] == 2'b11) begin
  anode <=4'b1000;
  cathode <= cat3;
 end

endmodule
